module moduleName (
    // IN
    input logic [2:0] alu_control,
    input logic [31:0] src1,
    input logic [31:0] scr2,
    // OUT
    output logic [31:0] alu_result,
    output logic zero
);

always_comb begin
    case (alu_control)
        3'b000 : alu_result = src1 + scr2;
        default: alu_result = 32'b0;
    endcase
end

assign zero = alu_result == 32'b0;
    
endmodule