module cpu (
    input logic clk,
    input logic rst,
    output logic [7:0] cnt
);
    
endmodule