/**
 *   HOLY_CLINT_AXI_LITE
 *
 *   Author : BRH
 *   Description : Pure Verilog wrapper for the Holy Core CLINT.
 *                 No SystemVerilog features. Ready for Vivado integration.
 */

module holy_clint_top #(
    parameter BASE_ADDR = 32'h0000_0000
)(
    input  wire                  clk,
    input  wire                  rst_n,

    // AXI Lite slave interface
    input  wire [31:0]           s_axi_awaddr,
    input  wire                  s_axi_awvalid,
    output wire                  s_axi_awready,
    input  wire [31:0]           s_axi_wdata,
    input  wire [3:0]            s_axi_wstrb,
    input  wire                  s_axi_wvalid,
    output wire                  s_axi_wready,
    output wire [1:0]            s_axi_bresp,
    output wire                  s_axi_bvalid,
    input  wire                  s_axi_bready,

    input  wire [31:0]           s_axi_araddr,
    input  wire                  s_axi_arvalid,
    output wire                  s_axi_arready,
    output wire [31:0]           s_axi_rdata,
    output wire [1:0]            s_axi_rresp,
    output wire                  s_axi_rvalid,
    input  wire                  s_axi_rready,

    // Interrupt outputs
    output wire                  timer_irq,
    output wire                  soft_irq
);

    // Instantiate stripped-down CLINT module
    holy_clint_wrapper #(
        .BASE_ADDR(BASE_ADDR)
    ) u_holy_clint_top (
        .clk(clk),
        .rst_n(rst_n),

        .s_axi_awaddr(s_axi_awaddr),
        .s_axi_awvalid(s_axi_awvalid),
        .s_axi_awready(s_axi_awready),
        .s_axi_wdata(s_axi_wdata),
        .s_axi_wstrb(s_axi_wstrb),
        .s_axi_wvalid(s_axi_wvalid),
        .s_axi_wready(s_axi_wready),
        .s_axi_bresp(s_axi_bresp),
        .s_axi_bvalid(s_axi_bvalid),
        .s_axi_bready(s_axi_bready),
        .s_axi_araddr(s_axi_araddr),
        .s_axi_arvalid(s_axi_arvalid),
        .s_axi_arready(s_axi_arready),
        .s_axi_rdata(s_axi_rdata),
        .s_axi_rresp(s_axi_rresp),
        .s_axi_rvalid(s_axi_rvalid),
        .s_axi_rready(s_axi_rready),

        .timer_irq(timer_irq),
        .soft_irq(soft_irq)
    );

endmodule
